library verilog;
use verilog.vl_types.all;
entity hazard_unit_sv_unit is
end hazard_unit_sv_unit;
